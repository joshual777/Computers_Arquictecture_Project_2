 module negador_1b (input logic a, output logic result );
										
assign result = ~a;

endmodule 